.OP 
Vc 1 0 5.008942 
C 6 8 1.033653u 
R1 1 2 1028.064358 
R2 3 2 2031.977037 
R3 2 5 3006.381471 
R4 5 0 4183.973331 
R5 6 5 3119.937426 
R6 4 7 2088.587447 
R7 7 8 1000.449867 
Gcs 6 3 2 5 0.007063 
Vprobe 0 4 0 
Hvs 5 8 Vprobe 8119.248145 
.END 
