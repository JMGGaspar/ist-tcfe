.OP 
**Voltage source ****************************************** 
Vcc vcc 0 12.000000 
Vin in 0 0 ac 1.0 sin(0 0.010000 1000.000000) 
Rin in in2 100.000000 

**coupling capacitor ****************************************** 
Ci in2 base  0.001000 

** bias circuit****************************************** 
Rb1 vcc base 80000.000000 
Rb2 base 0 20000.000000 

**gain stage ************************************* 
Q1 coll base emit BC547A 
Rc vcc coll 1000.000000 
Re emit 0 100.000000 

** bypass capacitor ************************************* 
Cb emit 0 0.001000 

**output stage ************************************* 
Q2 0 coll emit2 BC557A 
Rout emit2 vcc 100.000000 

**output coupling capacitor ************************************* 
Co emit2 out 0.000001 

**load ************************************* 
Rload out2 0 8.000000 
Vout out out2 0 

******************************************** 
.csparam Mu=2102.508000 

******************************************** 
.END 
