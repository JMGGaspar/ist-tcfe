.OP 
.param n={1/10.000000} 
**Voltage source ****************************************** 
Vc Ph 0  dc sin(0 230.000000 50.000000) 

**Transformer ****************************************** 
F1 Ph 0  E1  n 
E1 vac vacref Ph 0 n 

** Rectifier****************************************** 
DR1 vac 1 Default 
DR2 GND vac Default 
DR3 vacref 1 Default 
DR4 GND vacref Default 

**First regulation ************************************* 
C1 1 GND 15.000000u 
R1 1 GND 15.000000k 
R2 1 2 5.600000k 

**Final regulation**************************************** 
D1 2 3 Default 
D2 3 4 Default 
D3 4 5 Default 
D4 5 6 Default 
D5 6 7 Default 
D6 7 8 Default 
D7 8 9 Default 
D8 9 10 Default 
D9 10 11 Default 
D10 11 12 Default 
D11 12 13 Default 
D12 13 14 Default 
D13 14 15 Default 
D14 15 16 Default 
D15 16 17 Default 
D16 17 18 Default 
D17 18 19 Default 
D18 19 GND Default 

******************************************** 
.model Default D 
.csparam Mu=37.800000 

******************************************** 
.END 
